

architecture Behavioral of test_fixed_points is

begin


end Behavioral;
